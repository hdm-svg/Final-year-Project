`timescale 1ns/1ps
module linear_diffuse(
	input [63:0] x0,
	input [63:0] x1,
	input [63:0] x2,
	input [63:0] x3,
	input [63:0] x4,
	
	output [63:0] x0_o,
	output [63:0] x1_o,
	output [63:0] x2_o,
	output [63:0] x3_o,
	output [63:0] x4_o
);
	
	assign x0_o = x0 ^ {x0[18:0],x0[63:19]} ^ {x0[27:0],x0[63:28]};
	assign x1_o = x1 ^ {x1[60:0],x1[63:61]} ^ {x1[38:0],x1[63:39]};
	assign x2_o = x2 ^ {x2[0:0],x2[63:01]} ^ {x2[05:0],x2[63:06]};
	assign x3_o = x3 ^ {x3[9:0],x3[63:10]} ^ {x3[16:0],x3[63:17]};
	assign x4_o = x4 ^ {x4[6:0],x4[63:07]} ^ {x4[40:0],x4[63:41]};

//	assign x0_o = x0 ^ ((x0 >> 19) | ((x0 & (1<<19)-1) << (64-19))) ^ ((x0 >> 28) | ((x0 & (1<<28)-1) << (64-28)));
//	assign x1_o = x1 ^ ((x1 >> 61) | ((x1 & (1<<61)-1) << (64-61))) ^ ((x1 >> 39) | ((x1 & (1<<39)-1) << (64-39)));
//	assign x2_o = x2 ^ ((x2 >> 1)  | ((x2 & (1<<1)-1) << (64-1)))   ^ ((x2 >> 6)  | ((x2 & (1<<6)-1)  << (64-6)));
//	assign x3_o = x3 ^ ((x3 >> 10) | ((x3 & (1<<10)-1) << (64-10))) ^ ((x3 >> 17) | ((x3 & (1<<17)-1) << (64-17)));
//	assign x4_o = x4 ^ ((x4 >> 7)  | ((x4 & (1<<7)-1) << (64-7)))   ^ ((x4 >> 41) | ((x4 & (1<<41)-1) << (64-41)));

endmodule
